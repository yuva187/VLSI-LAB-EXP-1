module fs(a,b,bin,d,bout);
input a,b,bin;
output d,bout;



endmodule