module ha(a,b,sum,carry);
input a,b;
output sum,carry;

endmodule
